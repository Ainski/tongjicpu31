`timescale 1ns / 1ps
module sccomp_dataflow(
    input clk_in,
    input reset,
    output [31:0] NPCout,
    output [31:0] a,
    output [31:0] b,
    output [31:0] DMEMdata,
    output [31:0] imdt,
    output [25:0] index,
    output [31:0] inst,
    output [31:0] jextend,
    output [4:0] mux3out,
    output [31:0] npc,
    output [31:0] pc,
    output [31:0] rd,
    output [31:0] rdd,
    output [31:0] r,
    output [31:0] rs,
    output [31:0] rt,
    output [31:0] shamt,
    output [5:0] func,
    output [5:0] op,
    output [4:0] rdc,
    output [4:0] rsc,
    output [4:0] rtc,
    output [4:0] shamtT,
    output [3:0] aluc,
    output [3:0] jpc,
    output [15:0] imdtT,
    output [1:0] M1,
    output [1:0] M2,
    output [1:0] M3,
    output M4,
    output [1:0] M5,
    output Btype,
    output carry,
    output CS,
    output DM_R,
    output DM_W,
    output IM_R,
    output M6,
    output negative,
    output overflow,
    output RF_CLK,

    output RF_W,
    output su,
    output zero,
    output Ze,
    output [31:0] regfile0,regfile1,regfile2,regfile3,regfile4,regfile5,regfile6,regfile7,
    regfile8,regfile9,regfile10,regfile11,regfile12,regfile13,regfile14,regfile15,
    regfile16,regfile17,regfile18,regfile19,regfile20,regfile21,regfile22,regfile23,
    regfile24,regfile25,regfile26,regfile27,regfile28,regfile29,regfile30,regfile31
);
wire [31:0]pc_temp;
assign pc=pc_temp+32'h00400000;
assign RF_CLK = clk_in;
cpu sccpu(
        .clk(clk_in),
        .NPCout(NPCout),
        .a(a),
        .b(b),
        .DMEMdata(DMEMdata),
        .imdt(imdt),
        .index(index),
        .instr(inst),
        .jextend(jextend),
        .mux3out(mux3out),
        .npc(npc),
        .pc(pc_temp),
        .rd(rd),
        .rdd(rdd),
        .r(r),
        .rs(rs),
        .rt(rt),
        .shamt(shamt),
        .func(func),
        .op(op),
        .rdc(rdc),
        .rsc(rsc),
        .rtc(rtc),
        .shamtT(shamtT),
        .aluc(aluc),
        .jpc(jpc),
        .imdtT(imdtT),
        .M1(M1),
        .M2(M2),
        .M3(M3),
        .M4(M4),
        .M5(M5),
        .Btype(Btype),
        .carry(carry),
        .CS(CS),
        .DM_R(DM_R),
        .DM_W(DM_W),
        .IM_R(IM_R),
        .M6(M6),
        .negative(negative),
        .overflow(overflow),
        .RF_CLK(RF_CLK),
        .RF_W(RF_W),
        .reset(reset),
        .su(su),
        .zero(zero),
        .Ze(Ze),
        .regfile0(regfile0),
        .regfile1(regfile1),
        .regfile2(regfile2),
        .regfile3(regfile3),
        .regfile4(regfile4),
        .regfile5(regfile5),
        .regfile6(regfile6),
        .regfile7(regfile7),
        .regfile8(regfile8),
        .regfile9(regfile9),
        .regfile10(regfile10),
        .regfile11(regfile11),
        .regfile12(regfile12),
        .regfile13(regfile13),
        .regfile14(regfile14),
        .regfile15(regfile15),
        .regfile16(regfile16),
        .regfile17(regfile17),
        .regfile18(regfile18),
        .regfile19(regfile19),
        .regfile20(regfile20),
        .regfile21(regfile21),
        .regfile22(regfile22),
        .regfile23(regfile23),
        .regfile24(regfile24),
        .regfile25(regfile25),
        .regfile26(regfile26),
        .regfile27(regfile27),
        .regfile28(regfile28),
        .regfile29(regfile29),
        .regfile30(regfile30),
        .regfile31(regfile31)
);
DMEM dmem_inst(
    .CS(CS),
    .DM_R(DM_R),
    .DM_W(DM_W),
    .DMEMaddr(r),
    .DMEMdata(DMEMdata),
    .clk(clk_in),
    .rt(rt)
);
IMEM imem_inst(
    .IM_R(IM_R),
    .address(pc_temp),
    .func(func),
    .index(index),
    .instr(inst),
    .imdtT(imdtT),
    .op(op),
    .rdc(rdc),
    .rsc(rsc),
    .rtc(rtc),
    .shamtT(shamtT)
);


endmodule